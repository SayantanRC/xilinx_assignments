--------------------------------------------------------------------------------
-- Company: 
-- Engineer:
--
-- Create Date:   22:12:49 11/14/2018
-- Design Name:   
-- Module Name:   /home/sayantan/xilinx working dir/ass-1/full_adder_tb.vhd
-- Project Name:  ass-1
-- Target Device:  
-- Tool versions:  
-- Description:   
-- 
-- VHDL Test Bench Created by ISE for module: full_adder_using_half_adder
-- 
-- Dependencies:
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
-- Notes: 
-- This testbench has been automatically generated using types std_logic and
-- std_logic_vector for the ports of the unit under test.  Xilinx recommends
-- that these types always be used for the top-level I/O of a design in order
-- to guarantee that the testbench will bind correctly to the post-implementation 
-- simulation model.
--------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
 
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--USE ieee.numeric_std.ALL;
 
ENTITY full_adder_tb IS
END full_adder_tb;
 
ARCHITECTURE behavior OF full_adder_tb IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
    COMPONENT full_adder_using_half_adder
    PORT(
         A : IN  std_logic;
         B : IN  std_logic;
         Cin : IN  std_logic;
         S : OUT  std_logic;
         Cy : OUT  std_logic
        );
    END COMPONENT;
    

   --Inputs
   signal A : std_logic := '0';
   signal B : std_logic := '0';
   signal Cin : std_logic := '0';

 	--Outputs
   signal S : std_logic;
   signal Cy : std_logic;
   -- No clocks detected in port list. Replace <clock> below with 
   -- appropriate port name 
 
--   constant <clock>_period : time := 10 ns;
 
BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: full_adder_using_half_adder PORT MAP (
          A => A,
          B => B,
          Cin => Cin,
          S => S,
          Cy => Cy
        );

   -- Clock process definitions
--   <clock>_process :process
--   begin
--		<clock> <= '0';
--		wait for <clock>_period/2;
--		<clock> <= '1';
--		wait for <clock>_period/2;
--   end process;
 

   -- Stimulus process
   stim_proc: process
   begin		
      -- hold reset state for 100 ns.
--      wait for 100 ns;	

--      wait for <clock>_period*10;

      -- insert stimulus here 
		
		A <= '0';
		B <= '0';
		Cin <= '0';
		
		wait for 100 ns;	
		
		A <= '0';
		B <= '0';
		Cin <= '1';
		
		wait for 100 ns;	
		
		A <= '0';
		B <= '1';
		Cin <= '0';
		
		wait for 100 ns;	
		
		A <= '0';
		B <= '1';
		Cin <= '1';
		
		wait for 100 ns;	
		
		A <= '1';
		B <= '0';
		Cin <= '0';
		
		wait for 100 ns;	
		
		A <= '1';
		B <= '0';
		Cin <= '1';
		
		wait for 100 ns;	
		
		A <= '1';
		B <= '1';
		Cin <= '0';
		
		wait for 100 ns;	
		
		A <= '1';
		B <= '1';
		Cin <= '1';	

      wait;
   end process;

END;
